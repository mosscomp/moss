/*
Copyright 2020 The Moss Authors.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

`timescale 1ns / 1ps

module regfile (
    input clk,
    input write_ctrl,
    input [4:0] rs1,
    input [4:0] rs2,
    input [4:0] rd,
    input [63:0] data,
    output [63:0] rv1,
    output [63:0] rv2
);

  reg [63:0] registers[31:0];

  assign rv1 = registers[rs1];
  assign rv2 = registers[rs2];

  always @(posedge clk) begin
    if (write_ctrl) begin
      registers[rd] <= data;
    end
  end
endmodule
