/*
Copyright 2020 The Moss Authors.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

`timescale 1ns / 1ps

// ALU is passed a control signal and two arguments. It returns the result of
// the operation, which should be the same size as the arguments.
module alu (
    input [1:0] op,
    input [63:0] arg1,
    arg2,
    output reg [63:0] result
);

  // operations
  localparam OP_AND = 2'b00;
  localparam OP_OR = 2'b01;
  localparam OP_ADD = 2'b10;
  localparam OP_SUB = 2'b11;

  always @(op, arg1, arg2) begin
    case (op)
      OP_AND: begin
        result = arg1 & arg2;
      end
      OP_OR: begin
        result = arg1 | arg2;
      end
      OP_ADD: begin
        result = arg1 + arg2;
      end
      OP_SUB: begin
        result = arg1 - arg2;
      end
    endcase
  end
endmodule
